module not_32(S, A);
    input [31:0] A;
    output [31:0] S;

    not not1(S[0], A[0]);
    not not2(S[1], A[1]);
    not not3(S[2], A[2]);
    not not4(S[3], A[3]);
    not not5(S[4], A[4]);
    not not6(S[5], A[5]);
    not not7(S[6], A[6]);
    not not8(S[7], A[7]);
    not not9(S[8], A[8]);
    not not10(S[9], A[9]);
    not not11(S[10], A[10]);
    not not12(S[11], A[11]);
    not not13(S[12], A[12]);
    not not14(S[13], A[13]);
    not not15(S[14], A[14]);
    not not16(S[15], A[15]);
    not not17(S[16], A[16]);
    not not18(S[17], A[17]);
    not not19(S[18], A[18]);
    not not20(S[19], A[19]);
    not not21(S[20], A[20]);
    not not22(S[21], A[21]);
    not not23(S[22], A[22]);
    not not24(S[23], A[23]);
    not not25(S[24], A[24]);
    not not26(S[25], A[25]);
    not not27(S[26], A[26]);
    not not28(S[27], A[27]);
    not not29(S[28], A[28]);
    not not30(S[29], A[29]);
    not not31(S[30], A[30]);
    not not32(S[31], A[31]);

endmodule