module or_32(S, A, B);
    input [31:0] A, B;
    output [31:0] S;

    or A_B_or0(S[0], A[0], B[0]);
    or A_B_or1(S[1], A[1], B[1]);
    or A_B_or2(S[2], A[2], B[2]);
    or A_B_or3(S[3], A[3], B[3]);
    or A_B_or4(S[4], A[4], B[4]);
    or A_B_or5(S[5], A[5], B[5]);
    or A_B_or6(S[6], A[6], B[6]);
    or A_B_or7(S[7], A[7], B[7]);
    or A_B_or8(S[8], A[8], B[8]);
    or A_B_or9(S[9], A[9], B[9]);
    or A_B_or10(S[10], A[10], B[10]);
    or A_B_or11(S[11], A[11], B[11]);
    or A_B_or12(S[12], A[12], B[12]);
    or A_B_or13(S[13], A[13], B[13]);
    or A_B_or14(S[14], A[14], B[14]);
    or A_B_or15(S[15], A[15], B[15]);
    or A_B_or16(S[16], A[16], B[16]);
    or A_B_or17(S[17], A[17], B[17]);
    or A_B_or18(S[18], A[18], B[18]);
    or A_B_or19(S[19], A[19], B[19]);
    or A_B_or20(S[20], A[20], B[20]);
    or A_B_or21(S[21], A[21], B[21]);
    or A_B_or22(S[22], A[22], B[22]);
    or A_B_or23(S[23], A[23], B[23]);
    or A_B_or24(S[24], A[24], B[24]);
    or A_B_or25(S[25], A[25], B[25]);
    or A_B_or26(S[26], A[26], B[26]);
    or A_B_or27(S[27], A[27], B[27]);
    or A_B_or28(S[28], A[28], B[28]);
    or A_B_or29(S[29], A[29], B[29]);
    or A_B_or30(S[30], A[30], B[30]);
    or A_B_or31(S[31], A[31], B[31]);

endmodule